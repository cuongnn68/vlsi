module tb_memory();

endmodule