module top_level(
    clk,
    rst,
    en
);


endmodule